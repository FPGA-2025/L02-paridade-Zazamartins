module calcula_paridade (
  input [7:0] dado,
  output paridade
);

// implemente o seu código aqui

  assign paridade = ^dado;

endmodule
